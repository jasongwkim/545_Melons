`timescale 1ns / 1ps

module ti_mixer(
    input logic CLK,
    input logic [3:0] vol0, vol1, vol2, vol3,
    input logic [9:0] tone0, tone1, tone2
);

endmodule