//----------------------------------------------------------------------------
//  A-Z80 CPU Copyright (C) 2014,2016  Goran Devic, www.baltazarstudios.com
//
//  This program is free software; you can redistribute it and/or modify it
//  under the terms of the GNU General Public License as published by the Free
//  Software Foundation; either version 2 of the License, or (at your option)
//  any later version.
//
//  This program is distributed in the hope that it will be useful, but WITHOUT
//  ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
//  FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License for
//  more details.
//----------------------------------------------------------------------------
// Automatically generated by genref.py

// Module: control/decode_state.v
ctl_state_iy_set = 0;
ctl_state_ixiy_clr = 0;
ctl_state_ixiy_we = 0;
ctl_state_halt_set = 0;
ctl_state_tbl_clr = 0;
ctl_state_tbl_ed_set = 0;
ctl_state_tbl_cb_set = 0;
ctl_state_alu = 0;
ctl_repeat_we = 0;

// Module: control/interrupts.v
ctl_iff1_iff2 = 0;
ctl_iffx_we = 0;
ctl_iffx_bit = 0;
ctl_im_we = 0;
ctl_no_ints = 0;

// Module: control/ir.v
ctl_ir_we = 0;

// Module: control/memory_ifc.v
ctl_mRead = 0;
ctl_mWrite = 0;
ctl_iorw = 0;

// Module: alu/alu_control.v
ctl_shift_en = 0;
ctl_daa_oe = 0;
ctl_alu_op_low = 0;
ctl_cond_short = 0;
ctl_alu_core_hf = 0;
ctl_eval_cond = 0;
ctl_66_oe = 0;
ctl_pf_sel = 0;

// Module: alu/alu_select.v
ctl_alu_oe = 0;
ctl_alu_shift_oe = 0;
ctl_alu_op2_oe = 0;
ctl_alu_res_oe = 0;
ctl_alu_op1_oe = 0;
ctl_alu_bs_oe = 0;
ctl_alu_op1_sel_bus = 0;
ctl_alu_op1_sel_low = 0;
ctl_alu_op1_sel_zero = 0;
ctl_alu_op2_sel_zero = 0;
ctl_alu_op2_sel_bus = 0;
ctl_alu_op2_sel_lq = 0;
ctl_alu_sel_op2_neg = 0;
ctl_alu_sel_op2_high = 0;
ctl_alu_core_R = 0;
ctl_alu_core_V = 0;
ctl_alu_core_S = 0;

// Module: alu/alu_flags.v
ctl_flags_oe = 0;
ctl_flags_bus = 0;
ctl_flags_alu = 0;
ctl_flags_nf_set = 0;
ctl_flags_cf_set = 0;
ctl_flags_cf_cpl = 0;
ctl_flags_cf_we = 0;
ctl_flags_sz_we = 0;
ctl_flags_xy_we = 0;
ctl_flags_hf_we = 0;
ctl_flags_pf_we = 0;
ctl_flags_nf_we = 0;
ctl_flags_cf2_we = 0;
ctl_flags_hf_cpl = 0;
ctl_flags_use_cf2 = 0;
ctl_flags_hf2_we = 0;
ctl_flags_nf_clr = 0;
ctl_alu_zero_16bit = 0;
ctl_flags_cf2_sel_shift = 0;
ctl_flags_cf2_sel_daa = 0;

// Module: registers/reg_file.v
ctl_sw_4u = 0;
ctl_reg_in_hi = 0;
ctl_reg_in_lo = 0;
ctl_reg_out_lo = 0;
ctl_reg_out_hi = 0;

// Module: registers/reg_control.v
ctl_reg_exx = 0;
ctl_reg_ex_af = 0;
ctl_reg_ex_de_hl = 0;
ctl_reg_use_sp = 0;
ctl_reg_sel_pc = 0;
ctl_reg_sel_ir = 0;
ctl_reg_sel_wz = 0;
ctl_reg_gp_we = 0;
ctl_reg_not_pc = 0;
ctl_reg_sys_we_lo = 0;
ctl_reg_sys_we_hi = 0;
ctl_reg_sys_we = 0;
ctl_sw_4d = 0;
ctl_reg_gp_hilo = 0;
ctl_reg_gp_sel = 0;
ctl_reg_sys_hilo = 0;

// Module: bus/address_latch.v
ctl_inc_cy = 0;
ctl_inc_dec = 0;
ctl_al_we = 0;
ctl_inc_limit6 = 0;
ctl_bus_inc_oe = 0;
ctl_apin_mux = 0;
ctl_apin_mux2 = 0;

// Module: bus/bus_control.v
ctl_bus_ff_oe = 0;
ctl_bus_zero_oe = 0;

// Module: bus/bus_switch.v
ctl_sw_1u = 0;
ctl_sw_1d = 0;
ctl_sw_2u = 0;
ctl_sw_2d = 0;
ctl_sw_mask543_en = 0;

// Module: bus/data_pins.v
ctl_bus_db_we = 0;
ctl_bus_db_oe = 0;
